module Divisor(input wire [31:0] AFio, input wire [31:0] BFio, output wire [31:0] DivLoFio, output wire [31:0] DivHiFio);

assign DivLoFio = AFio;
assign DivHiFio = Bfio;

endmodule
